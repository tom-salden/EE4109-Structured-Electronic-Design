"Drive Capability CS-stage"
* C:\Users\tomsa\Documents\SturcturedElectronics2021\Chapter5\SLiCAP\cir\CSstageComponents.asc
R1 out 0 {R_L}
I1 0 N001 I value=0 dc=0 dcvar=0 noise=0
R2 N001 0 {R_s}
G1 out 0 N001 0 {g_m}
C1 N001 0 {c_gs+c_gb}
C2 out 0 {c_db}
C3 N001 out {c_dg}
R3 out 0 {1/g_o}
.param R_s=10G R_L=10k
.backanno
.end
