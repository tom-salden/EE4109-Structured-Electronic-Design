"Conclusion on the design process"
* E:\Universiteit\Master\7 Q2 - 2021\EE4109-Structured-Electronic-Design\cir\emptyCircuit.asc
V1 0 0 V
.backanno
.end
