"Assignment 3 - Noise analysis with flicker noise"
V1 N001 0 V value=0 dc=0 dcvar=0 noise=0
C1 N002 N001 {C_s}
XU1 N002 0 out NM18_noise ID={ID} IG={IG} W={W} L={L}
.param C_s=5p IG=0 ID=6.4m W=50u L=180n M=16
.lib SLiCAP.lib
.backanno
.end
