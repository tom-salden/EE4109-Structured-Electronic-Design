"Assignment 4 - Complementary-parallel CS output stage"
* E:\Universiteit\Master\7 Q2 - 2021\EE4109 - Structured Electronic Design\EE4109-Structured-Electronic-Design\cir\emptyCircuit.asc
V1 0 0 V
.backanno
.end
